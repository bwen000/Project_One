`timescale 1ns / 1ps

module find_min_delay_tb;
    reg [7:0] ascii_in;
    wire [7:0] ascii_out;
    
    toUpper uut(ascii_in, ascii_out);
    
    parameter DELAY = 26;
    
    initial begin
        $dumpfile("find_min_delay_tb.vcd");
        $dumpvars(0, find_min_delay_tb);
        
        $display("========================================");
        $display("Testing with inter-input delay = %0d ns", DELAY);
        $display("========================================\n");
        $display("Time(ns)\tInput\tOutput\tExpected\tResult");
        $display("--------\t-----\t------\t--------\t------");
        
        ascii_in = 8'd0;
        #30;
        
        ascii_in = 8'd40; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 40, (ascii_out==40)?"PASS":"FAIL");
        
        ascii_in = 8'd72; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 72, (ascii_out==72)?"PASS":"FAIL");
        
        ascii_in = 8'd183; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 183, (ascii_out==183)?"PASS":"FAIL");
        
        ascii_in = 8'd131; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 131, (ascii_out==131)?"PASS":"FAIL");
        
        ascii_in = 8'd124; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 124, (ascii_out==124)?"PASS":"FAIL");
        
        ascii_in = 8'd20; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 20, (ascii_out==20)?"PASS":"FAIL");
        
        ascii_in = 8'd235; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 235, (ascii_out==235)?"PASS":"FAIL");
        
        ascii_in = 8'd97; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 65, (ascii_out==65)?"PASS":"FAIL");
        
        ascii_in = 8'd65; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 65, (ascii_out==65)?"PASS":"FAIL");
        
        ascii_in = 8'd122; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 90, (ascii_out==90)?"PASS":"FAIL");
        
        ascii_in = 8'd71; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 71, (ascii_out==71)?"PASS":"FAIL");
        
        ascii_in = 8'd109; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 77, (ascii_out==77)?"PASS":"FAIL");
        
        ascii_in = 8'd146; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 146, (ascii_out==146)?"PASS":"FAIL");
        
        ascii_in = 8'd48; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 48, (ascii_out==48)?"PASS":"FAIL");
        
        ascii_in = 8'd207; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 207, (ascii_out==207)?"PASS":"FAIL");
        
        ascii_in = 8'd58; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 58, (ascii_out==58)?"PASS":"FAIL");
        
        ascii_in = 8'd123; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 123, (ascii_out==123)?"PASS":"FAIL");
        
        ascii_in = 8'd148; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 148, (ascii_out==148)?"PASS":"FAIL");
        
        ascii_in = 8'd127; #DELAY;
        $display("%0t\t\t%d\t%d\t%d\t\t%s", $time, ascii_in, ascii_out, 127, (ascii_out==127)?"PASS":"FAIL");
        
        #50;
        $display("\n========================================");
        $display("Test complete with delay = %0d ns", DELAY);
        $display("========================================");
        $finish;
    end
endmodule